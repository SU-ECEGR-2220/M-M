--------------------------------------------------------------------------------
--
-- LAB #4
--
--------------------------------------------------------------------------------

Library ieee;
Use ieee.std_logic_1164.all;
Use ieee.numeric_std.all;
Use ieee.std_logic_unsigned.all;

entity ALU is
	Port(	DataIn1: in std_logic_vector(31 downto 0);
		DataIn2: in std_logic_vector(31 downto 0);
		ALUCtrl: in std_logic_vector(4 downto 0);
		Zero: out std_logic;
		ALUResult: out std_logic_vector(31 downto 0) );
end entity ALU;

architecture ALU_Arch of ALU is
	-- ALU components	
	component adder_subtracter
		port(	datain_a: in std_logic_vector(31 downto 0);
			datain_b: in std_logic_vector(31 downto 0);
			add_sub: in std_logic;
			dataout: out std_logic_vector(31 downto 0);
			co: out std_logic);
	end component adder_subtracter;

	component shift_register
		port(	datain: in std_logic_vector(31 downto 0);
		   	dir: in std_logic;
			shamt:	in std_logic_vector(4 downto 0);
			dataout: out std_logic_vector(31 downto 0));
	end component shift_register;

begin
	-- Add ALU VHDL implementation here
	direction <= ALUCtrl(0) xor ALUCtrl(1);

	with ALUCtrl select
	copy <=		M1(31 downto 0) when "
			M2(31 downto 0) when "
			DataIn1 and DataIn2 when "
			DataIn1 or DataIn2 when"
			DataIn2(31 downto 0) when others;

	alu1: adder_subtracter port map(
	alu2: shift_register port map(

	ALUResult <= copy(31 downto 0);

	with copy select
	Zero <= '1' when "
		'0' when others;

end architecture ALU_Arch;


